* Flip-Flop
.param supply=1.0
.param t_r=10p
.param t_f=20p
.temp 70
.model pmos pmos VTH0='-0.3*supply' level=14
.model nmos nmos VTH0='0.3*supply' level=14
.global vdd gnd
.inc libs/cirs.cir
Vdd vdd 0 'supply'

* Voltage sources/ Signal sources
V1 en  0 PULSE 0 'supply' 0.1n 't_r' 't_f' 1n 5n
V2 nen 0 PULSE 'supply' 0 0.1n 't_r' 't_f' 1n 5n
V3 a 0 PULSE 0 'supply' 0.3n 't_r' 't_f' 1n 2n

* Buffer
X0 a q inv N=10
X1 q q_buf inv N=10

* master-slave ff active rising edge
X2 q_buf en nen q1 ff_r N=2
* master-slave ff active falling edge
X3 q_buf en nen q2 ff_f N=2

* * Output Buffers
* X4 q1 q1_bar inv N=10
* X5 q1_bar q1_buf inv N=10
* X6 q2 q2_bar inv N=10
* X7 q2_bar q2_buf inv N=10

C1 q1 0 10f
C2 q2 0 10f

.tran 20n
