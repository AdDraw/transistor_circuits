* XOR gate

.param supply=1.0
.param t_r=10p
.param t_f=20p
.temp 70
.model pmos pmos VTH0='-0.3*supply' level=14
.model nmos nmos VTH0='0.3*supply' level=14

.global vdd gnd
.inc libs/cirs.cir

* Vdd
Vdd vdd 0 'supply'
* input 1
Vin1 in1         0 PULSE 0 'supply' 0.1n 't_r' 't_f' 0.5n 1n
Vin2 in1_bar 0 PULSE 'supply' 0 0.1n 't_r' 't_f' 0.5n 1n
* input 2
Vin3 in2         0 PULSE 0 'supply' 0.1n 't_r' 't_f' 1n 2n
Vin4 in2_bar 0 PULSE 'supply' 0 0.1n 't_r' 't_f' 1n 2n

X1 in1 in2                               out1 xor2_nand        N=4
X2 in1 in2                               out2 xor2_nor           N=4
X3 in1 in1_bar in2  in2_bar out3 xor2_tran          N=4
X4 in1 in1_bar in2  in2_bar out4  xor2_tran_opt N=4

# load
C1 out1 0 10f
C2 out2 0 10f
C3 out3 0 10f
C4 out4 0 10f


.tran 10n
