* simple circuits as subckts

.subckt inv in out
  M1 out in vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 out in gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends inv

.subckt buf in out
  X0 in     in_bar inv N={N}
  X1 in_bar out    inv N={N}
.ends buf

.subckt nand2 in1 in2 out
  * PUN
  M1 out in1 vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 out in2 vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  * PDN
  M3 out in1 tmp gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M4 tmp in2 gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends nand2

.subckt nand3 in1 in2 in3 out
  * PUN
  M1 out in1 vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 out in2 vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M3 out in3 vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  * PDN
  M4 out  in1 tmp  gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M5 tmp  in2 tmp2 gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M6 tmp2 in3 gnd  gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends nand3

.subckt nor2 in1 in2 out
  * PUN
  M1 out in1 tmp vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 tmp in2 vdd vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  * PDN
  M3 out in1 gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M4 out in2 gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends nor2

.subckt nor3 in1 in2 in3 out
  * PUN
  M1 out  in1 tmp  vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 tmp  in2 tmp2 vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M3 tmp2 in3 vdd  vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  * PDN
  M4 out in1 gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M5 out in2 gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M6 out in3 gnd gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends nor3

.subckt xor2_nand A B Q
  X1 A B AB_bar nand2 N={N}
  X2 A AB_bar tmp1 nand2 N={N}
  X3 B AB_bar tmp2 nand2 N={N}
  X4 tmp1 tmp2 Q nand2 N={N}
.ends xor2_nand

.subckt xor2_nor A B Q
  X1 A B Q1 nor2 N={N}
  X2 A Q1 Q2 nor2 N={N}
  X3 B Q1 Q3 nor2 N={N}
  X4 Q3 Q2 Q4 nor2 N={N}
  X5 Q4 Q4 Q nor2 N={N}
.ends xor2_nor

.subckt xor2_tran A A_bar B B_bar Q
  * PUN
  M1 vdd  A     tmp0 vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 vdd  B     tmp0 vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M3 tmp0 A_bar Q    vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M4 tmp0 B_bar Q    vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  * PDN
  M5 Q    A     tmp1 gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M6 tmp1 B     gnd  gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M7 Q    A_bar tmp2 gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M8 tmp2 B_bar gnd  gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends xor2_tran

.subckt xor2_tran_opt A A_bar B B_bar Q
  * PUN
  M1 vdd  A     tmp1 vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 tmp1 B_bar Q    vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M3 vdd  A_bar tmp2 vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M4 tmp2 B     Q    vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  * PDN
  M5 Q    A     tmp3 gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M6 tmp3 B     gnd  gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M7 Q    A_bar tmp4 gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M8 tmp4 B_bar gnd  gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends xor2_tran_opt

.subckt tg in out en nen
  M1 in nen out vdd pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  M2 in en  out gnd nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends tg

.subckt d_latch d en nen q q_bar
  X0 d     q     en  nen tg  N={N}
  X1 q     q_bar         inv N={N}
  X2 q_bar q2            inv N={N}
  X3 q2    q     nen en  tg  N={N}
.ends d_latch


.subckt d_latch_alt1 d s en nen q q_bar
  X0 d     q     en  nen tg  N={N}
  X1 q     q_bar         inv N={N}
  X2 s q_bar q2          nand2 N={N}
  X3 q2    q     nen en  tg  N={N}
.ends d_latch_alt1

.subckt d_latch_alt3 d r en nen q q_bar
  X0 d     q     en  nen tg  N={N}
  X1 q     q_bar         inv N={N}
  X2 r q_bar q2          nor2 N={N}
  X3 q2    q     nen en  tg  N={N}
.ends d_latch_alt3

.subckt d_latch_alt2 d s en nen q q_bar
  X0 d  q  en  nen       tg N={N}
  X1 s q   q_bar         nand2 N={N}
  X2 q_bar q2            inv N={N}
  X3 q2    q     nen en  tg  N={N}
.ends d_latch_alt2

.subckt d_latch_alt4 d r en nen q q_bar
  X0 d  q  en  nen       tg N={N}
  X1 r q   q_bar         nor2 N={N}
  X2 q_bar q2            inv N={N}
  X3 q2    q     nen en  tg  N={N}
.ends d_latch_alt4

.subckt d_latch_with_async_reset_active_low d r en nen q q_bar
  X0 d r norq nand2       N={N}
  X1 norq q en nen tg     N={N}
  X2 q q_bar inv          N={N}
  X3 q_bar r norq2 nand2  N={N}
  X4 norq2 q nen en tg    N={N}
.ends d_latch_with_async_reset_active_low

.subckt d_latch_with_async_set_active_high d s en nen q q_bar
  X0 d s norq nor2        N={N}
  X1 norq q en nen tg     N={N}
  X2 q q_bar inv          N={N}
  X3 q_bar s norq2 nor2   N={N}
  X4 norq2 q nen en tg    N={N}
.ends d_latch_with_async_set_active_high

.subckt d_latch_async_ctrl_active_high d q q_bar en nen ctrl z
  * z- if 1 then SET, 0 - RESET
  Xmux0 d z ctrl mux0out mux21 N={N}
  Xtg0  mux0out q en nen tg N={N}
  Xinv0 q q_bar inv N={N}
  Xinv1 q_bar tmp inv N={N}
  Xmux1 tmp z ctrl mux1out mux21 N={N}
  Xtg1  mux1out q nen en tg N={N}
.ends

.subckt d_latch_async_ctrl_active_low d q q_bar en nen ctrl z
  * z- if 1 then SET, 0 - RESET
  Xmux0 z d ctrl mux0out mux21 N={N}
  Xtg0  mux0out q en nen tg N={N}
  Xinv0 q q_bar inv N={N}
  Xinv1 q_bar tmp inv N={N}
  Xmux1 z tmp ctrl mux1out mux21 N={N}
  Xtg1  mux1out q nen en tg N={N}
.ends

.subckt ff_r d en nen q
  * Master (active low)
  X_master d nen en mq mq_bar d_latch N={N}
  * Slave (active high)
  X_slave mq_bar en nen sq q d_latch N={N}
.ends ff_r

.subckt ffrls d s en nen q
  * Master (active low)
  X_master d s nen en mq mq_bar d_latch_alt1 N={N}
  * Slave (active high)
  X_slave mq_bar s en nen sq q d_latch_alt2 N={N}
.ends ffrls

.subckt ffrhr d r en nen q
  * Master (active low)
  X_master d r nen en mq mq_bar d_latch_alt3 N={N}
  * Slave (active high)
  X_slave mq_bar r en nen sq q d_latch_alt4 N={N}
.ends ffrhr

.subckt ff_f d en nen q
  * Master (active high)
  X_master d en nen mq mq_bar d_latch N={N}
  * Slave (active low)
  X_slave mq_bar nen en sq q d_latch N={N}
.ends ff_f

.subckt fffls d s en nen q
  * Master (active high)
  X_master d s en nen mq mq_bar d_latch_alt1 N={N}
  * Slave (active low)
  X_slave mq_bar s nen en sq q d_latch_alt2 N={N}
.ends fffls

.subckt fffhr d r en nen q
  * Master (active high)
  X_master d r en nen mq mq_bar d_latch_alt3 N={N}
  * Slave (active low)
  X_slave mq_bar r nen en sq q d_latch_alt4 N={N}
.ends fffls


.subckt MUX21 a b s q
  Xinv s s_bar inv N={N}
  X0   a q s_bar s tg N={N}
  X1   b q s s_bar tg N={N}
.ends


** XOR3 lib
.subckt serialp3 a b c top bot body
  Mpt top  a  tmp1 body pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  Mpm tmp1 b  tmp2 body pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  Mpb tmp2 c  bot  body pmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends

.subckt paralleln3 a b c top bot body
  Mpt top a bot body nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  Mpm top b bot body nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
  Mpb top c bot body nmos W=100n L=50n AD=0 AS=0 PD=0 PS=0 m={N}
.ends

.subckt XOR3 a b c q
  * INPUT INVERTERS
  Xinv0 a a_bar inv N={N}
  Xinv1 b b_bar inv N={N}
  Xinv2 c c_bar inv N={N}
  * PUN
  X0 a     b     c_bar vdd q vdd serialp3 N={N}
  X1 a     b_bar c     vdd q vdd serialp3 N={N}
  X2 a_bar b     c     vdd q vdd serialp3 N={N}
  X3 a_bar b_bar c_bar vdd q vdd serialp3 N={N}
  * PDN
  X4 a     b     c_bar q    tmp1 gnd paralleln3 N={N}
  X5 a     b_bar c     tmp1 tmp2 gnd paralleln3 N={N}
  X6 a_bar b     c     tmp2 tmp3 gnd paralleln3 N={N}
  X7 a_bar b_bar c_bar tmp3 gnd  gnd paralleln3 N={N}
.ends