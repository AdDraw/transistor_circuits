* simple NOR2 gate

.param supply=1.0
.temp 70
.model pmos pmos VTH0='-0.3*supply' level=14
.model nmos nmos VTH0='0.3*supply' level=14

.global vdd gnd
.inc libs/cirs.cir

* Vdd
Vdd vdd 0 'supply'
* input 1
Vin1 in1 0 PULSE 0 'supply' .45n 0.05n 0.05n 0.45n 1n
* input 2
Vin2 in2 0 PULSE 0 'supply' 1n 0.05n 0.05n 0.9n 2n

X1 in1 in2 out xor2 N=10
X2 out out_bar inv N=10

# load
C1 out 0 10f
C2 out_bar 0 10f

.tran 10n
