* Flip-Flop
.param supply=1.0
.param t_r=10p
.param t_f=20p
.temp 70
.model pmos pmos VTH0='-0.3*supply' level=14
.model nmos nmos VTH0='0.3*supply' level=14
.global vdd gnd
.inc libs/cirs.cir
Vdd vdd 0 'supply'

* Voltage sources/ Signal sources
V1 en  0 PULSE 0 'supply' 0.1n 't_r' 't_f' 1n 2n
V2 nen 0 PULSE 'supply' 0 0.1n 't_r' 't_f' 1n 2n
V3 a 0 PULSE 0 'supply' 0.3n 't_r' 't_f' 3n 6n
V4 sr 0 PULSE 0 'supply' 0n 't_r' 't_f' 15n 30n

* Buffer
X0 a q_buf buf N=10

* master-slave ff active rising edge
X2 q_buf en nen q1 ff_r N=2
* master-slave ff active rising edge, active low set
X3 q_buf sr en nen q2 ffrls N=2
* master-slave ff active rising edge, active high reset
X6 q_buf sr en nen q5 ffrhr N=2
* master-slave ff active falling edge
X4 q_buf en nen q3 ff_f N=2
* master-slave ff active falling edge, active low set
X5 q_buf sr en nen q4 fffls N=2
* master-slave ff active falling edge, active high reset
X7 q_buf sr en nen q6 fffhr N=2


C1 q1 0 10f
C2 q2 0 10f
C3 q3 0 10f
C4 q4 0 10f
C5 q5 0 10f
C6 q6  0 10f
.tran 30n
